`timescale 1ns/10ps
module t_sorting();
	reg [31:0] 	wire [31:0] 	sorting test(		#300
		$finish;
	end
endmodule
