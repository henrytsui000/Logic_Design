module checkbig(A, B, Q);
	input [31:0] A, B;
	output Q;
	wire [31:0] rev_B, bit, rev_xor, state;
	not not31(rev_B[31], B[31]);
	not not30(rev_B[30], B[30]);
	not not29(rev_B[29], B[29]);
	not not28(rev_B[28], B[28]);
	not not27(rev_B[27], B[27]);
	not not26(rev_B[26], B[26]);
	not not25(rev_B[25], B[25]);
	not not24(rev_B[24], B[24]);
	not not23(rev_B[23], B[23]);
	not not22(rev_B[22], B[22]);
	not not21(rev_B[21], B[21]);
	not not20(rev_B[20], B[20]);
	not not19(rev_B[19], B[19]);
	not not18(rev_B[18], B[18]);
	not not17(rev_B[17], B[17]);
	not not16(rev_B[16], B[16]);
	not not15(rev_B[15], B[15]);
	not not14(rev_B[14], B[14]);
	not not13(rev_B[13], B[13]);
	not not12(rev_B[12], B[12]);
	not not11(rev_B[11], B[11]);
	not not10(rev_B[10], B[10]);
	not not9(rev_B[9], B[9]);
	not not8(rev_B[8], B[8]);
	not not7(rev_B[7], B[7]);
	not not6(rev_B[6], B[6]);
	not not5(rev_B[5], B[5]);
	not not4(rev_B[4], B[4]);
	not not3(rev_B[3], B[3]);
	not not2(rev_B[2], B[2]);
	not not1(rev_B[1], B[1]);
	not not0(rev_B[0], B[0]);

	xor xor31(bit[31], A[31], B[31]);
	xor xor30(bit[30], A[30], B[30]);
	xor xor29(bit[29], A[29], B[29]);
	xor xor28(bit[28], A[28], B[28]);
	xor xor27(bit[27], A[27], B[27]);
	xor xor26(bit[26], A[26], B[26]);
	xor xor25(bit[25], A[25], B[25]);
	xor xor24(bit[24], A[24], B[24]);
	xor xor23(bit[23], A[23], B[23]);
	xor xor22(bit[22], A[22], B[22]);
	xor xor21(bit[21], A[21], B[21]);
	xor xor20(bit[20], A[20], B[20]);
	xor xor19(bit[19], A[19], B[19]);
	xor xor18(bit[18], A[18], B[18]);
	xor xor17(bit[17], A[17], B[17]);
	xor xor16(bit[16], A[16], B[16]);
	xor xor15(bit[15], A[15], B[15]);
	xor xor14(bit[14], A[14], B[14]);
	xor xor13(bit[13], A[13], B[13]);
	xor xor12(bit[12], A[12], B[12]);
	xor xor11(bit[11], A[11], B[11]);
	xor xor10(bit[10], A[10], B[10]);
	xor xor9(bit[9], A[9], B[9]);
	xor xor8(bit[8], A[8], B[8]);
	xor xor7(bit[7], A[7], B[7]);
	xor xor6(bit[6], A[6], B[6]);
	xor xor5(bit[5], A[5], B[5]);
	xor xor4(bit[4], A[4], B[4]);
	xor xor3(bit[3], A[3], B[3]);
	xor xor2(bit[2], A[2], B[2]);
	xor xor1(bit[1], A[1], B[1]);
	xor xor0(bit[0], A[0], B[0]);

	not not63(rev_xor[31], bit[31]);
	not not62(rev_xor[30], bit[30]);
	not not61(rev_xor[29], bit[29]);
	not not60(rev_xor[28], bit[28]);
	not not59(rev_xor[27], bit[27]);
	not not58(rev_xor[26], bit[26]);
	not not57(rev_xor[25], bit[25]);
	not not56(rev_xor[24], bit[24]);
	not not55(rev_xor[23], bit[23]);
	not not54(rev_xor[22], bit[22]);
	not not53(rev_xor[21], bit[21]);
	not not52(rev_xor[20], bit[20]);
	not not51(rev_xor[19], bit[19]);
	not not50(rev_xor[18], bit[18]);
	not not49(rev_xor[17], bit[17]);
	not not48(rev_xor[16], bit[16]);
	not not47(rev_xor[15], bit[15]);
	not not46(rev_xor[14], bit[14]);
	not not45(rev_xor[13], bit[13]);
	not not44(rev_xor[12], bit[12]);
	not not43(rev_xor[11], bit[11]);
	not not42(rev_xor[10], bit[10]);
	not not41(rev_xor[9], bit[9]);
	not not40(rev_xor[8], bit[8]);
	not not39(rev_xor[7], bit[7]);
	not not38(rev_xor[6], bit[6]);
	not not37(rev_xor[5], bit[5]);
	not not36(rev_xor[4], bit[4]);
	not not35(rev_xor[3], bit[3]);
	not not34(rev_xor[2], bit[2]);
	not not33(rev_xor[1], bit[1]);
	not not32(rev_xor[0], bit[0]);

	and and31(state[31], A[31], rev_B[31]);
	and and30(state[30], A[30], rev_B[30], rev_xor[31]);
	and and29(state[29], A[29], rev_B[29], rev_xor[31], rev_xor[30]);
	and and28(state[28], A[28], rev_B[28], rev_xor[31], rev_xor[30], rev_xor[29]);
	and and27(state[27], A[27], rev_B[27], rev_xor[31], rev_xor[30], rev_xor[29], rev_xor[28]);
	and and26(state[26], A[26], rev_B[26], rev_xor[31], rev_xor[30], rev_xor[29], rev_xor[28], rev_xor[27]);
	and and25(state[25], A[25], rev_B[25], rev_xor[31], rev_xor[30], rev_xor[29], rev_xor[28], rev_xor[27], rev_xor[26]);
	and and24(state[24], A[24], rev_B[24], rev_xor[31], rev_xor[30], rev_xor[29], rev_xor[28], rev_xor[27], rev_xor[26], rev_xor[25]);
	and and23(state[23], A[23], rev_B[23], rev_xor[31], rev_xor[30], rev_xor[29], rev_xor[28], rev_xor[27], rev_xor[26], rev_xor[25], rev_xor[24]);
	and and22(state[22], A[22], rev_B[22], rev_xor[31], rev_xor[30], rev_xor[29], rev_xor[28], rev_xor[27], rev_xor[26], rev_xor[25], rev_xor[24], rev_xor[23]);
	and and21(state[21], A[21], rev_B[21], rev_xor[31], rev_xor[30], rev_xor[29], rev_xor[28], rev_xor[27], rev_xor[26], rev_xor[25], rev_xor[24], rev_xor[23], rev_xor[22]);
	and and20(state[20], A[20], rev_B[20], rev_xor[31], rev_xor[30], rev_xor[29], rev_xor[28], rev_xor[27], rev_xor[26], rev_xor[25], rev_xor[24], rev_xor[23], rev_xor[22], rev_xor[21]);
	and and19(state[19], A[19], rev_B[19], rev_xor[31], rev_xor[30], rev_xor[29], rev_xor[28], rev_xor[27], rev_xor[26], rev_xor[25], rev_xor[24], rev_xor[23], rev_xor[22], rev_xor[21], rev_xor[20]);
	and and18(state[18], A[18], rev_B[18], rev_xor[31], rev_xor[30], rev_xor[29], rev_xor[28], rev_xor[27], rev_xor[26], rev_xor[25], rev_xor[24], rev_xor[23], rev_xor[22], rev_xor[21], rev_xor[20], rev_xor[19]);
	and and17(state[17], A[17], rev_B[17], rev_xor[31], rev_xor[30], rev_xor[29], rev_xor[28], rev_xor[27], rev_xor[26], rev_xor[25], rev_xor[24], rev_xor[23], rev_xor[22], rev_xor[21], rev_xor[20], rev_xor[19], rev_xor[18]);
	and and16(state[16], A[16], rev_B[16], rev_xor[31], rev_xor[30], rev_xor[29], rev_xor[28], rev_xor[27], rev_xor[26], rev_xor[25], rev_xor[24], rev_xor[23], rev_xor[22], rev_xor[21], rev_xor[20], rev_xor[19], rev_xor[18], rev_xor[17]);
	and and15(state[15], A[15], rev_B[15], rev_xor[31], rev_xor[30], rev_xor[29], rev_xor[28], rev_xor[27], rev_xor[26], rev_xor[25], rev_xor[24], rev_xor[23], rev_xor[22], rev_xor[21], rev_xor[20], rev_xor[19], rev_xor[18], rev_xor[17], rev_xor[16]);
	and and14(state[14], A[14], rev_B[14], rev_xor[31], rev_xor[30], rev_xor[29], rev_xor[28], rev_xor[27], rev_xor[26], rev_xor[25], rev_xor[24], rev_xor[23], rev_xor[22], rev_xor[21], rev_xor[20], rev_xor[19], rev_xor[18], rev_xor[17], rev_xor[16], rev_xor[15]);
	and and13(state[13], A[13], rev_B[13], rev_xor[31], rev_xor[30], rev_xor[29], rev_xor[28], rev_xor[27], rev_xor[26], rev_xor[25], rev_xor[24], rev_xor[23], rev_xor[22], rev_xor[21], rev_xor[20], rev_xor[19], rev_xor[18], rev_xor[17], rev_xor[16], rev_xor[15], rev_xor[14]);
	and and12(state[12], A[12], rev_B[12], rev_xor[31], rev_xor[30], rev_xor[29], rev_xor[28], rev_xor[27], rev_xor[26], rev_xor[25], rev_xor[24], rev_xor[23], rev_xor[22], rev_xor[21], rev_xor[20], rev_xor[19], rev_xor[18], rev_xor[17], rev_xor[16], rev_xor[15], rev_xor[14], rev_xor[13]);
	and and11(state[11], A[11], rev_B[11], rev_xor[31], rev_xor[30], rev_xor[29], rev_xor[28], rev_xor[27], rev_xor[26], rev_xor[25], rev_xor[24], rev_xor[23], rev_xor[22], rev_xor[21], rev_xor[20], rev_xor[19], rev_xor[18], rev_xor[17], rev_xor[16], rev_xor[15], rev_xor[14], rev_xor[13], rev_xor[12]);
	and and10(state[10], A[10], rev_B[10], rev_xor[31], rev_xor[30], rev_xor[29], rev_xor[28], rev_xor[27], rev_xor[26], rev_xor[25], rev_xor[24], rev_xor[23], rev_xor[22], rev_xor[21], rev_xor[20], rev_xor[19], rev_xor[18], rev_xor[17], rev_xor[16], rev_xor[15], rev_xor[14], rev_xor[13], rev_xor[12], rev_xor[11]);
	and and9(state[9], A[9], rev_B[9], rev_xor[31], rev_xor[30], rev_xor[29], rev_xor[28], rev_xor[27], rev_xor[26], rev_xor[25], rev_xor[24], rev_xor[23], rev_xor[22], rev_xor[21], rev_xor[20], rev_xor[19], rev_xor[18], rev_xor[17], rev_xor[16], rev_xor[15], rev_xor[14], rev_xor[13], rev_xor[12], rev_xor[11], rev_xor[10]);
	and and8(state[8], A[8], rev_B[8], rev_xor[31], rev_xor[30], rev_xor[29], rev_xor[28], rev_xor[27], rev_xor[26], rev_xor[25], rev_xor[24], rev_xor[23], rev_xor[22], rev_xor[21], rev_xor[20], rev_xor[19], rev_xor[18], rev_xor[17], rev_xor[16], rev_xor[15], rev_xor[14], rev_xor[13], rev_xor[12], rev_xor[11], rev_xor[10], rev_xor[9]);
	and and7(state[7], A[7], rev_B[7], rev_xor[31], rev_xor[30], rev_xor[29], rev_xor[28], rev_xor[27], rev_xor[26], rev_xor[25], rev_xor[24], rev_xor[23], rev_xor[22], rev_xor[21], rev_xor[20], rev_xor[19], rev_xor[18], rev_xor[17], rev_xor[16], rev_xor[15], rev_xor[14], rev_xor[13], rev_xor[12], rev_xor[11], rev_xor[10], rev_xor[9], rev_xor[8]);
	and and6(state[6], A[6], rev_B[6], rev_xor[31], rev_xor[30], rev_xor[29], rev_xor[28], rev_xor[27], rev_xor[26], rev_xor[25], rev_xor[24], rev_xor[23], rev_xor[22], rev_xor[21], rev_xor[20], rev_xor[19], rev_xor[18], rev_xor[17], rev_xor[16], rev_xor[15], rev_xor[14], rev_xor[13], rev_xor[12], rev_xor[11], rev_xor[10], rev_xor[9], rev_xor[8], rev_xor[7]);
	and and5(state[5], A[5], rev_B[5], rev_xor[31], rev_xor[30], rev_xor[29], rev_xor[28], rev_xor[27], rev_xor[26], rev_xor[25], rev_xor[24], rev_xor[23], rev_xor[22], rev_xor[21], rev_xor[20], rev_xor[19], rev_xor[18], rev_xor[17], rev_xor[16], rev_xor[15], rev_xor[14], rev_xor[13], rev_xor[12], rev_xor[11], rev_xor[10], rev_xor[9], rev_xor[8], rev_xor[7], rev_xor[6]);
	and and4(state[4], A[4], rev_B[4], rev_xor[31], rev_xor[30], rev_xor[29], rev_xor[28], rev_xor[27], rev_xor[26], rev_xor[25], rev_xor[24], rev_xor[23], rev_xor[22], rev_xor[21], rev_xor[20], rev_xor[19], rev_xor[18], rev_xor[17], rev_xor[16], rev_xor[15], rev_xor[14], rev_xor[13], rev_xor[12], rev_xor[11], rev_xor[10], rev_xor[9], rev_xor[8], rev_xor[7], rev_xor[6], rev_xor[5]);
	and and3(state[3], A[3], rev_B[3], rev_xor[31], rev_xor[30], rev_xor[29], rev_xor[28], rev_xor[27], rev_xor[26], rev_xor[25], rev_xor[24], rev_xor[23], rev_xor[22], rev_xor[21], rev_xor[20], rev_xor[19], rev_xor[18], rev_xor[17], rev_xor[16], rev_xor[15], rev_xor[14], rev_xor[13], rev_xor[12], rev_xor[11], rev_xor[10], rev_xor[9], rev_xor[8], rev_xor[7], rev_xor[6], rev_xor[5], rev_xor[4]);
	and and2(state[2], A[2], rev_B[2], rev_xor[31], rev_xor[30], rev_xor[29], rev_xor[28], rev_xor[27], rev_xor[26], rev_xor[25], rev_xor[24], rev_xor[23], rev_xor[22], rev_xor[21], rev_xor[20], rev_xor[19], rev_xor[18], rev_xor[17], rev_xor[16], rev_xor[15], rev_xor[14], rev_xor[13], rev_xor[12], rev_xor[11], rev_xor[10], rev_xor[9], rev_xor[8], rev_xor[7], rev_xor[6], rev_xor[5], rev_xor[4], rev_xor[3]);
	and and1(state[1], A[1], rev_B[1], rev_xor[31], rev_xor[30], rev_xor[29], rev_xor[28], rev_xor[27], rev_xor[26], rev_xor[25], rev_xor[24], rev_xor[23], rev_xor[22], rev_xor[21], rev_xor[20], rev_xor[19], rev_xor[18], rev_xor[17], rev_xor[16], rev_xor[15], rev_xor[14], rev_xor[13], rev_xor[12], rev_xor[11], rev_xor[10], rev_xor[9], rev_xor[8], rev_xor[7], rev_xor[6], rev_xor[5], rev_xor[4], rev_xor[3], rev_xor[2]);
	and and0(state[0], A[0], rev_B[0], rev_xor[31], rev_xor[30], rev_xor[29], rev_xor[28], rev_xor[27], rev_xor[26], rev_xor[25], rev_xor[24], rev_xor[23], rev_xor[22], rev_xor[21], rev_xor[20], rev_xor[19], rev_xor[18], rev_xor[17], rev_xor[16], rev_xor[15], rev_xor[14], rev_xor[13], rev_xor[12], rev_xor[11], rev_xor[10], rev_xor[9], rev_xor[8], rev_xor[7], rev_xor[6], rev_xor[5], rev_xor[4], rev_xor[3], rev_xor[2], rev_xor[1]);

	or ans(Q, state[31], state[30], state[29], state[28], state[27], state[26], state[25], state[24], state[23], state[22], state[21], state[20], state[19], state[18], state[17], state[16], state[15], state[14], state[13], state[12], state[11], state[10], state[9], state[8], state[7], state[6], state[5], state[4], state[3], state[2], state[1], state[0]);
endmodule