`include "checkbig.v"
`include "mux.v"
module sorting(	input [31:0] 	output [31:0] 
endmodule