module HW_5 #(parameter N = 8) (input [N-1:0]in,output wire [N-1:0]out);
assign out = in;
endmodule