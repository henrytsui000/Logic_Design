`include "adder.v"
module full_adder(A, B, Cin, sum, Cout);
	input[1023:0]A, B;
	input Cin;
	output [1023:0]sum;
	output Cout;

	wire W[1024:0];

	adder a1(A[0], B[0], Cin, sum[0], W[0]);
	adder a2(A[1], B[1], W[0], sum[1], W[1]);
	adder a3(A[2], B[2], W[1], sum[2], W[2]);
	adder a4(A[3], B[3], W[2], sum[3], W[3]);
	adder a5(A[4], B[4], W[3], sum[4], W[4]);
	adder a6(A[5], B[5], W[4], sum[5], W[5]);
	adder a7(A[6], B[6], W[5], sum[6], W[6]);
	adder a8(A[7], B[7], W[6], sum[7], W[7]);
	adder a9(A[8], B[8], W[7], sum[8], W[8]);
	adder a10(A[9], B[9], W[8], sum[9], W[9]);
	adder a11(A[10], B[10], W[9], sum[10], W[10]);
	adder a12(A[11], B[11], W[10], sum[11], W[11]);
	adder a13(A[12], B[12], W[11], sum[12], W[12]);
	adder a14(A[13], B[13], W[12], sum[13], W[13]);
	adder a15(A[14], B[14], W[13], sum[14], W[14]);
	adder a16(A[15], B[15], W[14], sum[15], W[15]);
	adder a17(A[16], B[16], W[15], sum[16], W[16]);
	adder a18(A[17], B[17], W[16], sum[17], W[17]);
	adder a19(A[18], B[18], W[17], sum[18], W[18]);
	adder a20(A[19], B[19], W[18], sum[19], W[19]);
	adder a21(A[20], B[20], W[19], sum[20], W[20]);
	adder a22(A[21], B[21], W[20], sum[21], W[21]);
	adder a23(A[22], B[22], W[21], sum[22], W[22]);
	adder a24(A[23], B[23], W[22], sum[23], W[23]);
	adder a25(A[24], B[24], W[23], sum[24], W[24]);
	adder a26(A[25], B[25], W[24], sum[25], W[25]);
	adder a27(A[26], B[26], W[25], sum[26], W[26]);
	adder a28(A[27], B[27], W[26], sum[27], W[27]);
	adder a29(A[28], B[28], W[27], sum[28], W[28]);
	adder a30(A[29], B[29], W[28], sum[29], W[29]);
	adder a31(A[30], B[30], W[29], sum[30], W[30]);
	adder a32(A[31], B[31], W[30], sum[31], W[31]);
	adder a33(A[32], B[32], W[31], sum[32], W[32]);
	adder a34(A[33], B[33], W[32], sum[33], W[33]);
	adder a35(A[34], B[34], W[33], sum[34], W[34]);
	adder a36(A[35], B[35], W[34], sum[35], W[35]);
	adder a37(A[36], B[36], W[35], sum[36], W[36]);
	adder a38(A[37], B[37], W[36], sum[37], W[37]);
	adder a39(A[38], B[38], W[37], sum[38], W[38]);
	adder a40(A[39], B[39], W[38], sum[39], W[39]);
	adder a41(A[40], B[40], W[39], sum[40], W[40]);
	adder a42(A[41], B[41], W[40], sum[41], W[41]);
	adder a43(A[42], B[42], W[41], sum[42], W[42]);
	adder a44(A[43], B[43], W[42], sum[43], W[43]);
	adder a45(A[44], B[44], W[43], sum[44], W[44]);
	adder a46(A[45], B[45], W[44], sum[45], W[45]);
	adder a47(A[46], B[46], W[45], sum[46], W[46]);
	adder a48(A[47], B[47], W[46], sum[47], W[47]);
	adder a49(A[48], B[48], W[47], sum[48], W[48]);
	adder a50(A[49], B[49], W[48], sum[49], W[49]);
	adder a51(A[50], B[50], W[49], sum[50], W[50]);
	adder a52(A[51], B[51], W[50], sum[51], W[51]);
	adder a53(A[52], B[52], W[51], sum[52], W[52]);
	adder a54(A[53], B[53], W[52], sum[53], W[53]);
	adder a55(A[54], B[54], W[53], sum[54], W[54]);
	adder a56(A[55], B[55], W[54], sum[55], W[55]);
	adder a57(A[56], B[56], W[55], sum[56], W[56]);
	adder a58(A[57], B[57], W[56], sum[57], W[57]);
	adder a59(A[58], B[58], W[57], sum[58], W[58]);
	adder a60(A[59], B[59], W[58], sum[59], W[59]);
	adder a61(A[60], B[60], W[59], sum[60], W[60]);
	adder a62(A[61], B[61], W[60], sum[61], W[61]);
	adder a63(A[62], B[62], W[61], sum[62], W[62]);
	adder a64(A[63], B[63], W[62], sum[63], W[63]);
	adder a65(A[64], B[64], W[63], sum[64], W[64]);
	adder a66(A[65], B[65], W[64], sum[65], W[65]);
	adder a67(A[66], B[66], W[65], sum[66], W[66]);
	adder a68(A[67], B[67], W[66], sum[67], W[67]);
	adder a69(A[68], B[68], W[67], sum[68], W[68]);
	adder a70(A[69], B[69], W[68], sum[69], W[69]);
	adder a71(A[70], B[70], W[69], sum[70], W[70]);
	adder a72(A[71], B[71], W[70], sum[71], W[71]);
	adder a73(A[72], B[72], W[71], sum[72], W[72]);
	adder a74(A[73], B[73], W[72], sum[73], W[73]);
	adder a75(A[74], B[74], W[73], sum[74], W[74]);
	adder a76(A[75], B[75], W[74], sum[75], W[75]);
	adder a77(A[76], B[76], W[75], sum[76], W[76]);
	adder a78(A[77], B[77], W[76], sum[77], W[77]);
	adder a79(A[78], B[78], W[77], sum[78], W[78]);
	adder a80(A[79], B[79], W[78], sum[79], W[79]);
	adder a81(A[80], B[80], W[79], sum[80], W[80]);
	adder a82(A[81], B[81], W[80], sum[81], W[81]);
	adder a83(A[82], B[82], W[81], sum[82], W[82]);
	adder a84(A[83], B[83], W[82], sum[83], W[83]);
	adder a85(A[84], B[84], W[83], sum[84], W[84]);
	adder a86(A[85], B[85], W[84], sum[85], W[85]);
	adder a87(A[86], B[86], W[85], sum[86], W[86]);
	adder a88(A[87], B[87], W[86], sum[87], W[87]);
	adder a89(A[88], B[88], W[87], sum[88], W[88]);
	adder a90(A[89], B[89], W[88], sum[89], W[89]);
	adder a91(A[90], B[90], W[89], sum[90], W[90]);
	adder a92(A[91], B[91], W[90], sum[91], W[91]);
	adder a93(A[92], B[92], W[91], sum[92], W[92]);
	adder a94(A[93], B[93], W[92], sum[93], W[93]);
	adder a95(A[94], B[94], W[93], sum[94], W[94]);
	adder a96(A[95], B[95], W[94], sum[95], W[95]);
	adder a97(A[96], B[96], W[95], sum[96], W[96]);
	adder a98(A[97], B[97], W[96], sum[97], W[97]);
	adder a99(A[98], B[98], W[97], sum[98], W[98]);
	adder a100(A[99], B[99], W[98], sum[99], W[99]);
	adder a101(A[100], B[100], W[99], sum[100], W[100]);
	adder a102(A[101], B[101], W[100], sum[101], W[101]);
	adder a103(A[102], B[102], W[101], sum[102], W[102]);
	adder a104(A[103], B[103], W[102], sum[103], W[103]);
	adder a105(A[104], B[104], W[103], sum[104], W[104]);
	adder a106(A[105], B[105], W[104], sum[105], W[105]);
	adder a107(A[106], B[106], W[105], sum[106], W[106]);
	adder a108(A[107], B[107], W[106], sum[107], W[107]);
	adder a109(A[108], B[108], W[107], sum[108], W[108]);
	adder a110(A[109], B[109], W[108], sum[109], W[109]);
	adder a111(A[110], B[110], W[109], sum[110], W[110]);
	adder a112(A[111], B[111], W[110], sum[111], W[111]);
	adder a113(A[112], B[112], W[111], sum[112], W[112]);
	adder a114(A[113], B[113], W[112], sum[113], W[113]);
	adder a115(A[114], B[114], W[113], sum[114], W[114]);
	adder a116(A[115], B[115], W[114], sum[115], W[115]);
	adder a117(A[116], B[116], W[115], sum[116], W[116]);
	adder a118(A[117], B[117], W[116], sum[117], W[117]);
	adder a119(A[118], B[118], W[117], sum[118], W[118]);
	adder a120(A[119], B[119], W[118], sum[119], W[119]);
	adder a121(A[120], B[120], W[119], sum[120], W[120]);
	adder a122(A[121], B[121], W[120], sum[121], W[121]);
	adder a123(A[122], B[122], W[121], sum[122], W[122]);
	adder a124(A[123], B[123], W[122], sum[123], W[123]);
	adder a125(A[124], B[124], W[123], sum[124], W[124]);
	adder a126(A[125], B[125], W[124], sum[125], W[125]);
	adder a127(A[126], B[126], W[125], sum[126], W[126]);
	adder a128(A[127], B[127], W[126], sum[127], W[127]);
	adder a129(A[128], B[128], W[127], sum[128], W[128]);
	adder a130(A[129], B[129], W[128], sum[129], W[129]);
	adder a131(A[130], B[130], W[129], sum[130], W[130]);
	adder a132(A[131], B[131], W[130], sum[131], W[131]);
	adder a133(A[132], B[132], W[131], sum[132], W[132]);
	adder a134(A[133], B[133], W[132], sum[133], W[133]);
	adder a135(A[134], B[134], W[133], sum[134], W[134]);
	adder a136(A[135], B[135], W[134], sum[135], W[135]);
	adder a137(A[136], B[136], W[135], sum[136], W[136]);
	adder a138(A[137], B[137], W[136], sum[137], W[137]);
	adder a139(A[138], B[138], W[137], sum[138], W[138]);
	adder a140(A[139], B[139], W[138], sum[139], W[139]);
	adder a141(A[140], B[140], W[139], sum[140], W[140]);
	adder a142(A[141], B[141], W[140], sum[141], W[141]);
	adder a143(A[142], B[142], W[141], sum[142], W[142]);
	adder a144(A[143], B[143], W[142], sum[143], W[143]);
	adder a145(A[144], B[144], W[143], sum[144], W[144]);
	adder a146(A[145], B[145], W[144], sum[145], W[145]);
	adder a147(A[146], B[146], W[145], sum[146], W[146]);
	adder a148(A[147], B[147], W[146], sum[147], W[147]);
	adder a149(A[148], B[148], W[147], sum[148], W[148]);
	adder a150(A[149], B[149], W[148], sum[149], W[149]);
	adder a151(A[150], B[150], W[149], sum[150], W[150]);
	adder a152(A[151], B[151], W[150], sum[151], W[151]);
	adder a153(A[152], B[152], W[151], sum[152], W[152]);
	adder a154(A[153], B[153], W[152], sum[153], W[153]);
	adder a155(A[154], B[154], W[153], sum[154], W[154]);
	adder a156(A[155], B[155], W[154], sum[155], W[155]);
	adder a157(A[156], B[156], W[155], sum[156], W[156]);
	adder a158(A[157], B[157], W[156], sum[157], W[157]);
	adder a159(A[158], B[158], W[157], sum[158], W[158]);
	adder a160(A[159], B[159], W[158], sum[159], W[159]);
	adder a161(A[160], B[160], W[159], sum[160], W[160]);
	adder a162(A[161], B[161], W[160], sum[161], W[161]);
	adder a163(A[162], B[162], W[161], sum[162], W[162]);
	adder a164(A[163], B[163], W[162], sum[163], W[163]);
	adder a165(A[164], B[164], W[163], sum[164], W[164]);
	adder a166(A[165], B[165], W[164], sum[165], W[165]);
	adder a167(A[166], B[166], W[165], sum[166], W[166]);
	adder a168(A[167], B[167], W[166], sum[167], W[167]);
	adder a169(A[168], B[168], W[167], sum[168], W[168]);
	adder a170(A[169], B[169], W[168], sum[169], W[169]);
	adder a171(A[170], B[170], W[169], sum[170], W[170]);
	adder a172(A[171], B[171], W[170], sum[171], W[171]);
	adder a173(A[172], B[172], W[171], sum[172], W[172]);
	adder a174(A[173], B[173], W[172], sum[173], W[173]);
	adder a175(A[174], B[174], W[173], sum[174], W[174]);
	adder a176(A[175], B[175], W[174], sum[175], W[175]);
	adder a177(A[176], B[176], W[175], sum[176], W[176]);
	adder a178(A[177], B[177], W[176], sum[177], W[177]);
	adder a179(A[178], B[178], W[177], sum[178], W[178]);
	adder a180(A[179], B[179], W[178], sum[179], W[179]);
	adder a181(A[180], B[180], W[179], sum[180], W[180]);
	adder a182(A[181], B[181], W[180], sum[181], W[181]);
	adder a183(A[182], B[182], W[181], sum[182], W[182]);
	adder a184(A[183], B[183], W[182], sum[183], W[183]);
	adder a185(A[184], B[184], W[183], sum[184], W[184]);
	adder a186(A[185], B[185], W[184], sum[185], W[185]);
	adder a187(A[186], B[186], W[185], sum[186], W[186]);
	adder a188(A[187], B[187], W[186], sum[187], W[187]);
	adder a189(A[188], B[188], W[187], sum[188], W[188]);
	adder a190(A[189], B[189], W[188], sum[189], W[189]);
	adder a191(A[190], B[190], W[189], sum[190], W[190]);
	adder a192(A[191], B[191], W[190], sum[191], W[191]);
	adder a193(A[192], B[192], W[191], sum[192], W[192]);
	adder a194(A[193], B[193], W[192], sum[193], W[193]);
	adder a195(A[194], B[194], W[193], sum[194], W[194]);
	adder a196(A[195], B[195], W[194], sum[195], W[195]);
	adder a197(A[196], B[196], W[195], sum[196], W[196]);
	adder a198(A[197], B[197], W[196], sum[197], W[197]);
	adder a199(A[198], B[198], W[197], sum[198], W[198]);
	adder a200(A[199], B[199], W[198], sum[199], W[199]);
	adder a201(A[200], B[200], W[199], sum[200], W[200]);
	adder a202(A[201], B[201], W[200], sum[201], W[201]);
	adder a203(A[202], B[202], W[201], sum[202], W[202]);
	adder a204(A[203], B[203], W[202], sum[203], W[203]);
	adder a205(A[204], B[204], W[203], sum[204], W[204]);
	adder a206(A[205], B[205], W[204], sum[205], W[205]);
	adder a207(A[206], B[206], W[205], sum[206], W[206]);
	adder a208(A[207], B[207], W[206], sum[207], W[207]);
	adder a209(A[208], B[208], W[207], sum[208], W[208]);
	adder a210(A[209], B[209], W[208], sum[209], W[209]);
	adder a211(A[210], B[210], W[209], sum[210], W[210]);
	adder a212(A[211], B[211], W[210], sum[211], W[211]);
	adder a213(A[212], B[212], W[211], sum[212], W[212]);
	adder a214(A[213], B[213], W[212], sum[213], W[213]);
	adder a215(A[214], B[214], W[213], sum[214], W[214]);
	adder a216(A[215], B[215], W[214], sum[215], W[215]);
	adder a217(A[216], B[216], W[215], sum[216], W[216]);
	adder a218(A[217], B[217], W[216], sum[217], W[217]);
	adder a219(A[218], B[218], W[217], sum[218], W[218]);
	adder a220(A[219], B[219], W[218], sum[219], W[219]);
	adder a221(A[220], B[220], W[219], sum[220], W[220]);
	adder a222(A[221], B[221], W[220], sum[221], W[221]);
	adder a223(A[222], B[222], W[221], sum[222], W[222]);
	adder a224(A[223], B[223], W[222], sum[223], W[223]);
	adder a225(A[224], B[224], W[223], sum[224], W[224]);
	adder a226(A[225], B[225], W[224], sum[225], W[225]);
	adder a227(A[226], B[226], W[225], sum[226], W[226]);
	adder a228(A[227], B[227], W[226], sum[227], W[227]);
	adder a229(A[228], B[228], W[227], sum[228], W[228]);
	adder a230(A[229], B[229], W[228], sum[229], W[229]);
	adder a231(A[230], B[230], W[229], sum[230], W[230]);
	adder a232(A[231], B[231], W[230], sum[231], W[231]);
	adder a233(A[232], B[232], W[231], sum[232], W[232]);
	adder a234(A[233], B[233], W[232], sum[233], W[233]);
	adder a235(A[234], B[234], W[233], sum[234], W[234]);
	adder a236(A[235], B[235], W[234], sum[235], W[235]);
	adder a237(A[236], B[236], W[235], sum[236], W[236]);
	adder a238(A[237], B[237], W[236], sum[237], W[237]);
	adder a239(A[238], B[238], W[237], sum[238], W[238]);
	adder a240(A[239], B[239], W[238], sum[239], W[239]);
	adder a241(A[240], B[240], W[239], sum[240], W[240]);
	adder a242(A[241], B[241], W[240], sum[241], W[241]);
	adder a243(A[242], B[242], W[241], sum[242], W[242]);
	adder a244(A[243], B[243], W[242], sum[243], W[243]);
	adder a245(A[244], B[244], W[243], sum[244], W[244]);
	adder a246(A[245], B[245], W[244], sum[245], W[245]);
	adder a247(A[246], B[246], W[245], sum[246], W[246]);
	adder a248(A[247], B[247], W[246], sum[247], W[247]);
	adder a249(A[248], B[248], W[247], sum[248], W[248]);
	adder a250(A[249], B[249], W[248], sum[249], W[249]);
	adder a251(A[250], B[250], W[249], sum[250], W[250]);
	adder a252(A[251], B[251], W[250], sum[251], W[251]);
	adder a253(A[252], B[252], W[251], sum[252], W[252]);
	adder a254(A[253], B[253], W[252], sum[253], W[253]);
	adder a255(A[254], B[254], W[253], sum[254], W[254]);
	adder a256(A[255], B[255], W[254], sum[255], W[255]);
	adder a257(A[256], B[256], W[255], sum[256], W[256]);
	adder a258(A[257], B[257], W[256], sum[257], W[257]);
	adder a259(A[258], B[258], W[257], sum[258], W[258]);
	adder a260(A[259], B[259], W[258], sum[259], W[259]);
	adder a261(A[260], B[260], W[259], sum[260], W[260]);
	adder a262(A[261], B[261], W[260], sum[261], W[261]);
	adder a263(A[262], B[262], W[261], sum[262], W[262]);
	adder a264(A[263], B[263], W[262], sum[263], W[263]);
	adder a265(A[264], B[264], W[263], sum[264], W[264]);
	adder a266(A[265], B[265], W[264], sum[265], W[265]);
	adder a267(A[266], B[266], W[265], sum[266], W[266]);
	adder a268(A[267], B[267], W[266], sum[267], W[267]);
	adder a269(A[268], B[268], W[267], sum[268], W[268]);
	adder a270(A[269], B[269], W[268], sum[269], W[269]);
	adder a271(A[270], B[270], W[269], sum[270], W[270]);
	adder a272(A[271], B[271], W[270], sum[271], W[271]);
	adder a273(A[272], B[272], W[271], sum[272], W[272]);
	adder a274(A[273], B[273], W[272], sum[273], W[273]);
	adder a275(A[274], B[274], W[273], sum[274], W[274]);
	adder a276(A[275], B[275], W[274], sum[275], W[275]);
	adder a277(A[276], B[276], W[275], sum[276], W[276]);
	adder a278(A[277], B[277], W[276], sum[277], W[277]);
	adder a279(A[278], B[278], W[277], sum[278], W[278]);
	adder a280(A[279], B[279], W[278], sum[279], W[279]);
	adder a281(A[280], B[280], W[279], sum[280], W[280]);
	adder a282(A[281], B[281], W[280], sum[281], W[281]);
	adder a283(A[282], B[282], W[281], sum[282], W[282]);
	adder a284(A[283], B[283], W[282], sum[283], W[283]);
	adder a285(A[284], B[284], W[283], sum[284], W[284]);
	adder a286(A[285], B[285], W[284], sum[285], W[285]);
	adder a287(A[286], B[286], W[285], sum[286], W[286]);
	adder a288(A[287], B[287], W[286], sum[287], W[287]);
	adder a289(A[288], B[288], W[287], sum[288], W[288]);
	adder a290(A[289], B[289], W[288], sum[289], W[289]);
	adder a291(A[290], B[290], W[289], sum[290], W[290]);
	adder a292(A[291], B[291], W[290], sum[291], W[291]);
	adder a293(A[292], B[292], W[291], sum[292], W[292]);
	adder a294(A[293], B[293], W[292], sum[293], W[293]);
	adder a295(A[294], B[294], W[293], sum[294], W[294]);
	adder a296(A[295], B[295], W[294], sum[295], W[295]);
	adder a297(A[296], B[296], W[295], sum[296], W[296]);
	adder a298(A[297], B[297], W[296], sum[297], W[297]);
	adder a299(A[298], B[298], W[297], sum[298], W[298]);
	adder a300(A[299], B[299], W[298], sum[299], W[299]);
	adder a301(A[300], B[300], W[299], sum[300], W[300]);
	adder a302(A[301], B[301], W[300], sum[301], W[301]);
	adder a303(A[302], B[302], W[301], sum[302], W[302]);
	adder a304(A[303], B[303], W[302], sum[303], W[303]);
	adder a305(A[304], B[304], W[303], sum[304], W[304]);
	adder a306(A[305], B[305], W[304], sum[305], W[305]);
	adder a307(A[306], B[306], W[305], sum[306], W[306]);
	adder a308(A[307], B[307], W[306], sum[307], W[307]);
	adder a309(A[308], B[308], W[307], sum[308], W[308]);
	adder a310(A[309], B[309], W[308], sum[309], W[309]);
	adder a311(A[310], B[310], W[309], sum[310], W[310]);
	adder a312(A[311], B[311], W[310], sum[311], W[311]);
	adder a313(A[312], B[312], W[311], sum[312], W[312]);
	adder a314(A[313], B[313], W[312], sum[313], W[313]);
	adder a315(A[314], B[314], W[313], sum[314], W[314]);
	adder a316(A[315], B[315], W[314], sum[315], W[315]);
	adder a317(A[316], B[316], W[315], sum[316], W[316]);
	adder a318(A[317], B[317], W[316], sum[317], W[317]);
	adder a319(A[318], B[318], W[317], sum[318], W[318]);
	adder a320(A[319], B[319], W[318], sum[319], W[319]);
	adder a321(A[320], B[320], W[319], sum[320], W[320]);
	adder a322(A[321], B[321], W[320], sum[321], W[321]);
	adder a323(A[322], B[322], W[321], sum[322], W[322]);
	adder a324(A[323], B[323], W[322], sum[323], W[323]);
	adder a325(A[324], B[324], W[323], sum[324], W[324]);
	adder a326(A[325], B[325], W[324], sum[325], W[325]);
	adder a327(A[326], B[326], W[325], sum[326], W[326]);
	adder a328(A[327], B[327], W[326], sum[327], W[327]);
	adder a329(A[328], B[328], W[327], sum[328], W[328]);
	adder a330(A[329], B[329], W[328], sum[329], W[329]);
	adder a331(A[330], B[330], W[329], sum[330], W[330]);
	adder a332(A[331], B[331], W[330], sum[331], W[331]);
	adder a333(A[332], B[332], W[331], sum[332], W[332]);
	adder a334(A[333], B[333], W[332], sum[333], W[333]);
	adder a335(A[334], B[334], W[333], sum[334], W[334]);
	adder a336(A[335], B[335], W[334], sum[335], W[335]);
	adder a337(A[336], B[336], W[335], sum[336], W[336]);
	adder a338(A[337], B[337], W[336], sum[337], W[337]);
	adder a339(A[338], B[338], W[337], sum[338], W[338]);
	adder a340(A[339], B[339], W[338], sum[339], W[339]);
	adder a341(A[340], B[340], W[339], sum[340], W[340]);
	adder a342(A[341], B[341], W[340], sum[341], W[341]);
	adder a343(A[342], B[342], W[341], sum[342], W[342]);
	adder a344(A[343], B[343], W[342], sum[343], W[343]);
	adder a345(A[344], B[344], W[343], sum[344], W[344]);
	adder a346(A[345], B[345], W[344], sum[345], W[345]);
	adder a347(A[346], B[346], W[345], sum[346], W[346]);
	adder a348(A[347], B[347], W[346], sum[347], W[347]);
	adder a349(A[348], B[348], W[347], sum[348], W[348]);
	adder a350(A[349], B[349], W[348], sum[349], W[349]);
	adder a351(A[350], B[350], W[349], sum[350], W[350]);
	adder a352(A[351], B[351], W[350], sum[351], W[351]);
	adder a353(A[352], B[352], W[351], sum[352], W[352]);
	adder a354(A[353], B[353], W[352], sum[353], W[353]);
	adder a355(A[354], B[354], W[353], sum[354], W[354]);
	adder a356(A[355], B[355], W[354], sum[355], W[355]);
	adder a357(A[356], B[356], W[355], sum[356], W[356]);
	adder a358(A[357], B[357], W[356], sum[357], W[357]);
	adder a359(A[358], B[358], W[357], sum[358], W[358]);
	adder a360(A[359], B[359], W[358], sum[359], W[359]);
	adder a361(A[360], B[360], W[359], sum[360], W[360]);
	adder a362(A[361], B[361], W[360], sum[361], W[361]);
	adder a363(A[362], B[362], W[361], sum[362], W[362]);
	adder a364(A[363], B[363], W[362], sum[363], W[363]);
	adder a365(A[364], B[364], W[363], sum[364], W[364]);
	adder a366(A[365], B[365], W[364], sum[365], W[365]);
	adder a367(A[366], B[366], W[365], sum[366], W[366]);
	adder a368(A[367], B[367], W[366], sum[367], W[367]);
	adder a369(A[368], B[368], W[367], sum[368], W[368]);
	adder a370(A[369], B[369], W[368], sum[369], W[369]);
	adder a371(A[370], B[370], W[369], sum[370], W[370]);
	adder a372(A[371], B[371], W[370], sum[371], W[371]);
	adder a373(A[372], B[372], W[371], sum[372], W[372]);
	adder a374(A[373], B[373], W[372], sum[373], W[373]);
	adder a375(A[374], B[374], W[373], sum[374], W[374]);
	adder a376(A[375], B[375], W[374], sum[375], W[375]);
	adder a377(A[376], B[376], W[375], sum[376], W[376]);
	adder a378(A[377], B[377], W[376], sum[377], W[377]);
	adder a379(A[378], B[378], W[377], sum[378], W[378]);
	adder a380(A[379], B[379], W[378], sum[379], W[379]);
	adder a381(A[380], B[380], W[379], sum[380], W[380]);
	adder a382(A[381], B[381], W[380], sum[381], W[381]);
	adder a383(A[382], B[382], W[381], sum[382], W[382]);
	adder a384(A[383], B[383], W[382], sum[383], W[383]);
	adder a385(A[384], B[384], W[383], sum[384], W[384]);
	adder a386(A[385], B[385], W[384], sum[385], W[385]);
	adder a387(A[386], B[386], W[385], sum[386], W[386]);
	adder a388(A[387], B[387], W[386], sum[387], W[387]);
	adder a389(A[388], B[388], W[387], sum[388], W[388]);
	adder a390(A[389], B[389], W[388], sum[389], W[389]);
	adder a391(A[390], B[390], W[389], sum[390], W[390]);
	adder a392(A[391], B[391], W[390], sum[391], W[391]);
	adder a393(A[392], B[392], W[391], sum[392], W[392]);
	adder a394(A[393], B[393], W[392], sum[393], W[393]);
	adder a395(A[394], B[394], W[393], sum[394], W[394]);
	adder a396(A[395], B[395], W[394], sum[395], W[395]);
	adder a397(A[396], B[396], W[395], sum[396], W[396]);
	adder a398(A[397], B[397], W[396], sum[397], W[397]);
	adder a399(A[398], B[398], W[397], sum[398], W[398]);
	adder a400(A[399], B[399], W[398], sum[399], W[399]);
	adder a401(A[400], B[400], W[399], sum[400], W[400]);
	adder a402(A[401], B[401], W[400], sum[401], W[401]);
	adder a403(A[402], B[402], W[401], sum[402], W[402]);
	adder a404(A[403], B[403], W[402], sum[403], W[403]);
	adder a405(A[404], B[404], W[403], sum[404], W[404]);
	adder a406(A[405], B[405], W[404], sum[405], W[405]);
	adder a407(A[406], B[406], W[405], sum[406], W[406]);
	adder a408(A[407], B[407], W[406], sum[407], W[407]);
	adder a409(A[408], B[408], W[407], sum[408], W[408]);
	adder a410(A[409], B[409], W[408], sum[409], W[409]);
	adder a411(A[410], B[410], W[409], sum[410], W[410]);
	adder a412(A[411], B[411], W[410], sum[411], W[411]);
	adder a413(A[412], B[412], W[411], sum[412], W[412]);
	adder a414(A[413], B[413], W[412], sum[413], W[413]);
	adder a415(A[414], B[414], W[413], sum[414], W[414]);
	adder a416(A[415], B[415], W[414], sum[415], W[415]);
	adder a417(A[416], B[416], W[415], sum[416], W[416]);
	adder a418(A[417], B[417], W[416], sum[417], W[417]);
	adder a419(A[418], B[418], W[417], sum[418], W[418]);
	adder a420(A[419], B[419], W[418], sum[419], W[419]);
	adder a421(A[420], B[420], W[419], sum[420], W[420]);
	adder a422(A[421], B[421], W[420], sum[421], W[421]);
	adder a423(A[422], B[422], W[421], sum[422], W[422]);
	adder a424(A[423], B[423], W[422], sum[423], W[423]);
	adder a425(A[424], B[424], W[423], sum[424], W[424]);
	adder a426(A[425], B[425], W[424], sum[425], W[425]);
	adder a427(A[426], B[426], W[425], sum[426], W[426]);
	adder a428(A[427], B[427], W[426], sum[427], W[427]);
	adder a429(A[428], B[428], W[427], sum[428], W[428]);
	adder a430(A[429], B[429], W[428], sum[429], W[429]);
	adder a431(A[430], B[430], W[429], sum[430], W[430]);
	adder a432(A[431], B[431], W[430], sum[431], W[431]);
	adder a433(A[432], B[432], W[431], sum[432], W[432]);
	adder a434(A[433], B[433], W[432], sum[433], W[433]);
	adder a435(A[434], B[434], W[433], sum[434], W[434]);
	adder a436(A[435], B[435], W[434], sum[435], W[435]);
	adder a437(A[436], B[436], W[435], sum[436], W[436]);
	adder a438(A[437], B[437], W[436], sum[437], W[437]);
	adder a439(A[438], B[438], W[437], sum[438], W[438]);
	adder a440(A[439], B[439], W[438], sum[439], W[439]);
	adder a441(A[440], B[440], W[439], sum[440], W[440]);
	adder a442(A[441], B[441], W[440], sum[441], W[441]);
	adder a443(A[442], B[442], W[441], sum[442], W[442]);
	adder a444(A[443], B[443], W[442], sum[443], W[443]);
	adder a445(A[444], B[444], W[443], sum[444], W[444]);
	adder a446(A[445], B[445], W[444], sum[445], W[445]);
	adder a447(A[446], B[446], W[445], sum[446], W[446]);
	adder a448(A[447], B[447], W[446], sum[447], W[447]);
	adder a449(A[448], B[448], W[447], sum[448], W[448]);
	adder a450(A[449], B[449], W[448], sum[449], W[449]);
	adder a451(A[450], B[450], W[449], sum[450], W[450]);
	adder a452(A[451], B[451], W[450], sum[451], W[451]);
	adder a453(A[452], B[452], W[451], sum[452], W[452]);
	adder a454(A[453], B[453], W[452], sum[453], W[453]);
	adder a455(A[454], B[454], W[453], sum[454], W[454]);
	adder a456(A[455], B[455], W[454], sum[455], W[455]);
	adder a457(A[456], B[456], W[455], sum[456], W[456]);
	adder a458(A[457], B[457], W[456], sum[457], W[457]);
	adder a459(A[458], B[458], W[457], sum[458], W[458]);
	adder a460(A[459], B[459], W[458], sum[459], W[459]);
	adder a461(A[460], B[460], W[459], sum[460], W[460]);
	adder a462(A[461], B[461], W[460], sum[461], W[461]);
	adder a463(A[462], B[462], W[461], sum[462], W[462]);
	adder a464(A[463], B[463], W[462], sum[463], W[463]);
	adder a465(A[464], B[464], W[463], sum[464], W[464]);
	adder a466(A[465], B[465], W[464], sum[465], W[465]);
	adder a467(A[466], B[466], W[465], sum[466], W[466]);
	adder a468(A[467], B[467], W[466], sum[467], W[467]);
	adder a469(A[468], B[468], W[467], sum[468], W[468]);
	adder a470(A[469], B[469], W[468], sum[469], W[469]);
	adder a471(A[470], B[470], W[469], sum[470], W[470]);
	adder a472(A[471], B[471], W[470], sum[471], W[471]);
	adder a473(A[472], B[472], W[471], sum[472], W[472]);
	adder a474(A[473], B[473], W[472], sum[473], W[473]);
	adder a475(A[474], B[474], W[473], sum[474], W[474]);
	adder a476(A[475], B[475], W[474], sum[475], W[475]);
	adder a477(A[476], B[476], W[475], sum[476], W[476]);
	adder a478(A[477], B[477], W[476], sum[477], W[477]);
	adder a479(A[478], B[478], W[477], sum[478], W[478]);
	adder a480(A[479], B[479], W[478], sum[479], W[479]);
	adder a481(A[480], B[480], W[479], sum[480], W[480]);
	adder a482(A[481], B[481], W[480], sum[481], W[481]);
	adder a483(A[482], B[482], W[481], sum[482], W[482]);
	adder a484(A[483], B[483], W[482], sum[483], W[483]);
	adder a485(A[484], B[484], W[483], sum[484], W[484]);
	adder a486(A[485], B[485], W[484], sum[485], W[485]);
	adder a487(A[486], B[486], W[485], sum[486], W[486]);
	adder a488(A[487], B[487], W[486], sum[487], W[487]);
	adder a489(A[488], B[488], W[487], sum[488], W[488]);
	adder a490(A[489], B[489], W[488], sum[489], W[489]);
	adder a491(A[490], B[490], W[489], sum[490], W[490]);
	adder a492(A[491], B[491], W[490], sum[491], W[491]);
	adder a493(A[492], B[492], W[491], sum[492], W[492]);
	adder a494(A[493], B[493], W[492], sum[493], W[493]);
	adder a495(A[494], B[494], W[493], sum[494], W[494]);
	adder a496(A[495], B[495], W[494], sum[495], W[495]);
	adder a497(A[496], B[496], W[495], sum[496], W[496]);
	adder a498(A[497], B[497], W[496], sum[497], W[497]);
	adder a499(A[498], B[498], W[497], sum[498], W[498]);
	adder a500(A[499], B[499], W[498], sum[499], W[499]);
	adder a501(A[500], B[500], W[499], sum[500], W[500]);
	adder a502(A[501], B[501], W[500], sum[501], W[501]);
	adder a503(A[502], B[502], W[501], sum[502], W[502]);
	adder a504(A[503], B[503], W[502], sum[503], W[503]);
	adder a505(A[504], B[504], W[503], sum[504], W[504]);
	adder a506(A[505], B[505], W[504], sum[505], W[505]);
	adder a507(A[506], B[506], W[505], sum[506], W[506]);
	adder a508(A[507], B[507], W[506], sum[507], W[507]);
	adder a509(A[508], B[508], W[507], sum[508], W[508]);
	adder a510(A[509], B[509], W[508], sum[509], W[509]);
	adder a511(A[510], B[510], W[509], sum[510], W[510]);
	adder a512(A[511], B[511], W[510], sum[511], W[511]);
	adder a513(A[512], B[512], W[511], sum[512], W[512]);
	adder a514(A[513], B[513], W[512], sum[513], W[513]);
	adder a515(A[514], B[514], W[513], sum[514], W[514]);
	adder a516(A[515], B[515], W[514], sum[515], W[515]);
	adder a517(A[516], B[516], W[515], sum[516], W[516]);
	adder a518(A[517], B[517], W[516], sum[517], W[517]);
	adder a519(A[518], B[518], W[517], sum[518], W[518]);
	adder a520(A[519], B[519], W[518], sum[519], W[519]);
	adder a521(A[520], B[520], W[519], sum[520], W[520]);
	adder a522(A[521], B[521], W[520], sum[521], W[521]);
	adder a523(A[522], B[522], W[521], sum[522], W[522]);
	adder a524(A[523], B[523], W[522], sum[523], W[523]);
	adder a525(A[524], B[524], W[523], sum[524], W[524]);
	adder a526(A[525], B[525], W[524], sum[525], W[525]);
	adder a527(A[526], B[526], W[525], sum[526], W[526]);
	adder a528(A[527], B[527], W[526], sum[527], W[527]);
	adder a529(A[528], B[528], W[527], sum[528], W[528]);
	adder a530(A[529], B[529], W[528], sum[529], W[529]);
	adder a531(A[530], B[530], W[529], sum[530], W[530]);
	adder a532(A[531], B[531], W[530], sum[531], W[531]);
	adder a533(A[532], B[532], W[531], sum[532], W[532]);
	adder a534(A[533], B[533], W[532], sum[533], W[533]);
	adder a535(A[534], B[534], W[533], sum[534], W[534]);
	adder a536(A[535], B[535], W[534], sum[535], W[535]);
	adder a537(A[536], B[536], W[535], sum[536], W[536]);
	adder a538(A[537], B[537], W[536], sum[537], W[537]);
	adder a539(A[538], B[538], W[537], sum[538], W[538]);
	adder a540(A[539], B[539], W[538], sum[539], W[539]);
	adder a541(A[540], B[540], W[539], sum[540], W[540]);
	adder a542(A[541], B[541], W[540], sum[541], W[541]);
	adder a543(A[542], B[542], W[541], sum[542], W[542]);
	adder a544(A[543], B[543], W[542], sum[543], W[543]);
	adder a545(A[544], B[544], W[543], sum[544], W[544]);
	adder a546(A[545], B[545], W[544], sum[545], W[545]);
	adder a547(A[546], B[546], W[545], sum[546], W[546]);
	adder a548(A[547], B[547], W[546], sum[547], W[547]);
	adder a549(A[548], B[548], W[547], sum[548], W[548]);
	adder a550(A[549], B[549], W[548], sum[549], W[549]);
	adder a551(A[550], B[550], W[549], sum[550], W[550]);
	adder a552(A[551], B[551], W[550], sum[551], W[551]);
	adder a553(A[552], B[552], W[551], sum[552], W[552]);
	adder a554(A[553], B[553], W[552], sum[553], W[553]);
	adder a555(A[554], B[554], W[553], sum[554], W[554]);
	adder a556(A[555], B[555], W[554], sum[555], W[555]);
	adder a557(A[556], B[556], W[555], sum[556], W[556]);
	adder a558(A[557], B[557], W[556], sum[557], W[557]);
	adder a559(A[558], B[558], W[557], sum[558], W[558]);
	adder a560(A[559], B[559], W[558], sum[559], W[559]);
	adder a561(A[560], B[560], W[559], sum[560], W[560]);
	adder a562(A[561], B[561], W[560], sum[561], W[561]);
	adder a563(A[562], B[562], W[561], sum[562], W[562]);
	adder a564(A[563], B[563], W[562], sum[563], W[563]);
	adder a565(A[564], B[564], W[563], sum[564], W[564]);
	adder a566(A[565], B[565], W[564], sum[565], W[565]);
	adder a567(A[566], B[566], W[565], sum[566], W[566]);
	adder a568(A[567], B[567], W[566], sum[567], W[567]);
	adder a569(A[568], B[568], W[567], sum[568], W[568]);
	adder a570(A[569], B[569], W[568], sum[569], W[569]);
	adder a571(A[570], B[570], W[569], sum[570], W[570]);
	adder a572(A[571], B[571], W[570], sum[571], W[571]);
	adder a573(A[572], B[572], W[571], sum[572], W[572]);
	adder a574(A[573], B[573], W[572], sum[573], W[573]);
	adder a575(A[574], B[574], W[573], sum[574], W[574]);
	adder a576(A[575], B[575], W[574], sum[575], W[575]);
	adder a577(A[576], B[576], W[575], sum[576], W[576]);
	adder a578(A[577], B[577], W[576], sum[577], W[577]);
	adder a579(A[578], B[578], W[577], sum[578], W[578]);
	adder a580(A[579], B[579], W[578], sum[579], W[579]);
	adder a581(A[580], B[580], W[579], sum[580], W[580]);
	adder a582(A[581], B[581], W[580], sum[581], W[581]);
	adder a583(A[582], B[582], W[581], sum[582], W[582]);
	adder a584(A[583], B[583], W[582], sum[583], W[583]);
	adder a585(A[584], B[584], W[583], sum[584], W[584]);
	adder a586(A[585], B[585], W[584], sum[585], W[585]);
	adder a587(A[586], B[586], W[585], sum[586], W[586]);
	adder a588(A[587], B[587], W[586], sum[587], W[587]);
	adder a589(A[588], B[588], W[587], sum[588], W[588]);
	adder a590(A[589], B[589], W[588], sum[589], W[589]);
	adder a591(A[590], B[590], W[589], sum[590], W[590]);
	adder a592(A[591], B[591], W[590], sum[591], W[591]);
	adder a593(A[592], B[592], W[591], sum[592], W[592]);
	adder a594(A[593], B[593], W[592], sum[593], W[593]);
	adder a595(A[594], B[594], W[593], sum[594], W[594]);
	adder a596(A[595], B[595], W[594], sum[595], W[595]);
	adder a597(A[596], B[596], W[595], sum[596], W[596]);
	adder a598(A[597], B[597], W[596], sum[597], W[597]);
	adder a599(A[598], B[598], W[597], sum[598], W[598]);
	adder a600(A[599], B[599], W[598], sum[599], W[599]);
	adder a601(A[600], B[600], W[599], sum[600], W[600]);
	adder a602(A[601], B[601], W[600], sum[601], W[601]);
	adder a603(A[602], B[602], W[601], sum[602], W[602]);
	adder a604(A[603], B[603], W[602], sum[603], W[603]);
	adder a605(A[604], B[604], W[603], sum[604], W[604]);
	adder a606(A[605], B[605], W[604], sum[605], W[605]);
	adder a607(A[606], B[606], W[605], sum[606], W[606]);
	adder a608(A[607], B[607], W[606], sum[607], W[607]);
	adder a609(A[608], B[608], W[607], sum[608], W[608]);
	adder a610(A[609], B[609], W[608], sum[609], W[609]);
	adder a611(A[610], B[610], W[609], sum[610], W[610]);
	adder a612(A[611], B[611], W[610], sum[611], W[611]);
	adder a613(A[612], B[612], W[611], sum[612], W[612]);
	adder a614(A[613], B[613], W[612], sum[613], W[613]);
	adder a615(A[614], B[614], W[613], sum[614], W[614]);
	adder a616(A[615], B[615], W[614], sum[615], W[615]);
	adder a617(A[616], B[616], W[615], sum[616], W[616]);
	adder a618(A[617], B[617], W[616], sum[617], W[617]);
	adder a619(A[618], B[618], W[617], sum[618], W[618]);
	adder a620(A[619], B[619], W[618], sum[619], W[619]);
	adder a621(A[620], B[620], W[619], sum[620], W[620]);
	adder a622(A[621], B[621], W[620], sum[621], W[621]);
	adder a623(A[622], B[622], W[621], sum[622], W[622]);
	adder a624(A[623], B[623], W[622], sum[623], W[623]);
	adder a625(A[624], B[624], W[623], sum[624], W[624]);
	adder a626(A[625], B[625], W[624], sum[625], W[625]);
	adder a627(A[626], B[626], W[625], sum[626], W[626]);
	adder a628(A[627], B[627], W[626], sum[627], W[627]);
	adder a629(A[628], B[628], W[627], sum[628], W[628]);
	adder a630(A[629], B[629], W[628], sum[629], W[629]);
	adder a631(A[630], B[630], W[629], sum[630], W[630]);
	adder a632(A[631], B[631], W[630], sum[631], W[631]);
	adder a633(A[632], B[632], W[631], sum[632], W[632]);
	adder a634(A[633], B[633], W[632], sum[633], W[633]);
	adder a635(A[634], B[634], W[633], sum[634], W[634]);
	adder a636(A[635], B[635], W[634], sum[635], W[635]);
	adder a637(A[636], B[636], W[635], sum[636], W[636]);
	adder a638(A[637], B[637], W[636], sum[637], W[637]);
	adder a639(A[638], B[638], W[637], sum[638], W[638]);
	adder a640(A[639], B[639], W[638], sum[639], W[639]);
	adder a641(A[640], B[640], W[639], sum[640], W[640]);
	adder a642(A[641], B[641], W[640], sum[641], W[641]);
	adder a643(A[642], B[642], W[641], sum[642], W[642]);
	adder a644(A[643], B[643], W[642], sum[643], W[643]);
	adder a645(A[644], B[644], W[643], sum[644], W[644]);
	adder a646(A[645], B[645], W[644], sum[645], W[645]);
	adder a647(A[646], B[646], W[645], sum[646], W[646]);
	adder a648(A[647], B[647], W[646], sum[647], W[647]);
	adder a649(A[648], B[648], W[647], sum[648], W[648]);
	adder a650(A[649], B[649], W[648], sum[649], W[649]);
	adder a651(A[650], B[650], W[649], sum[650], W[650]);
	adder a652(A[651], B[651], W[650], sum[651], W[651]);
	adder a653(A[652], B[652], W[651], sum[652], W[652]);
	adder a654(A[653], B[653], W[652], sum[653], W[653]);
	adder a655(A[654], B[654], W[653], sum[654], W[654]);
	adder a656(A[655], B[655], W[654], sum[655], W[655]);
	adder a657(A[656], B[656], W[655], sum[656], W[656]);
	adder a658(A[657], B[657], W[656], sum[657], W[657]);
	adder a659(A[658], B[658], W[657], sum[658], W[658]);
	adder a660(A[659], B[659], W[658], sum[659], W[659]);
	adder a661(A[660], B[660], W[659], sum[660], W[660]);
	adder a662(A[661], B[661], W[660], sum[661], W[661]);
	adder a663(A[662], B[662], W[661], sum[662], W[662]);
	adder a664(A[663], B[663], W[662], sum[663], W[663]);
	adder a665(A[664], B[664], W[663], sum[664], W[664]);
	adder a666(A[665], B[665], W[664], sum[665], W[665]);
	adder a667(A[666], B[666], W[665], sum[666], W[666]);
	adder a668(A[667], B[667], W[666], sum[667], W[667]);
	adder a669(A[668], B[668], W[667], sum[668], W[668]);
	adder a670(A[669], B[669], W[668], sum[669], W[669]);
	adder a671(A[670], B[670], W[669], sum[670], W[670]);
	adder a672(A[671], B[671], W[670], sum[671], W[671]);
	adder a673(A[672], B[672], W[671], sum[672], W[672]);
	adder a674(A[673], B[673], W[672], sum[673], W[673]);
	adder a675(A[674], B[674], W[673], sum[674], W[674]);
	adder a676(A[675], B[675], W[674], sum[675], W[675]);
	adder a677(A[676], B[676], W[675], sum[676], W[676]);
	adder a678(A[677], B[677], W[676], sum[677], W[677]);
	adder a679(A[678], B[678], W[677], sum[678], W[678]);
	adder a680(A[679], B[679], W[678], sum[679], W[679]);
	adder a681(A[680], B[680], W[679], sum[680], W[680]);
	adder a682(A[681], B[681], W[680], sum[681], W[681]);
	adder a683(A[682], B[682], W[681], sum[682], W[682]);
	adder a684(A[683], B[683], W[682], sum[683], W[683]);
	adder a685(A[684], B[684], W[683], sum[684], W[684]);
	adder a686(A[685], B[685], W[684], sum[685], W[685]);
	adder a687(A[686], B[686], W[685], sum[686], W[686]);
	adder a688(A[687], B[687], W[686], sum[687], W[687]);
	adder a689(A[688], B[688], W[687], sum[688], W[688]);
	adder a690(A[689], B[689], W[688], sum[689], W[689]);
	adder a691(A[690], B[690], W[689], sum[690], W[690]);
	adder a692(A[691], B[691], W[690], sum[691], W[691]);
	adder a693(A[692], B[692], W[691], sum[692], W[692]);
	adder a694(A[693], B[693], W[692], sum[693], W[693]);
	adder a695(A[694], B[694], W[693], sum[694], W[694]);
	adder a696(A[695], B[695], W[694], sum[695], W[695]);
	adder a697(A[696], B[696], W[695], sum[696], W[696]);
	adder a698(A[697], B[697], W[696], sum[697], W[697]);
	adder a699(A[698], B[698], W[697], sum[698], W[698]);
	adder a700(A[699], B[699], W[698], sum[699], W[699]);
	adder a701(A[700], B[700], W[699], sum[700], W[700]);
	adder a702(A[701], B[701], W[700], sum[701], W[701]);
	adder a703(A[702], B[702], W[701], sum[702], W[702]);
	adder a704(A[703], B[703], W[702], sum[703], W[703]);
	adder a705(A[704], B[704], W[703], sum[704], W[704]);
	adder a706(A[705], B[705], W[704], sum[705], W[705]);
	adder a707(A[706], B[706], W[705], sum[706], W[706]);
	adder a708(A[707], B[707], W[706], sum[707], W[707]);
	adder a709(A[708], B[708], W[707], sum[708], W[708]);
	adder a710(A[709], B[709], W[708], sum[709], W[709]);
	adder a711(A[710], B[710], W[709], sum[710], W[710]);
	adder a712(A[711], B[711], W[710], sum[711], W[711]);
	adder a713(A[712], B[712], W[711], sum[712], W[712]);
	adder a714(A[713], B[713], W[712], sum[713], W[713]);
	adder a715(A[714], B[714], W[713], sum[714], W[714]);
	adder a716(A[715], B[715], W[714], sum[715], W[715]);
	adder a717(A[716], B[716], W[715], sum[716], W[716]);
	adder a718(A[717], B[717], W[716], sum[717], W[717]);
	adder a719(A[718], B[718], W[717], sum[718], W[718]);
	adder a720(A[719], B[719], W[718], sum[719], W[719]);
	adder a721(A[720], B[720], W[719], sum[720], W[720]);
	adder a722(A[721], B[721], W[720], sum[721], W[721]);
	adder a723(A[722], B[722], W[721], sum[722], W[722]);
	adder a724(A[723], B[723], W[722], sum[723], W[723]);
	adder a725(A[724], B[724], W[723], sum[724], W[724]);
	adder a726(A[725], B[725], W[724], sum[725], W[725]);
	adder a727(A[726], B[726], W[725], sum[726], W[726]);
	adder a728(A[727], B[727], W[726], sum[727], W[727]);
	adder a729(A[728], B[728], W[727], sum[728], W[728]);
	adder a730(A[729], B[729], W[728], sum[729], W[729]);
	adder a731(A[730], B[730], W[729], sum[730], W[730]);
	adder a732(A[731], B[731], W[730], sum[731], W[731]);
	adder a733(A[732], B[732], W[731], sum[732], W[732]);
	adder a734(A[733], B[733], W[732], sum[733], W[733]);
	adder a735(A[734], B[734], W[733], sum[734], W[734]);
	adder a736(A[735], B[735], W[734], sum[735], W[735]);
	adder a737(A[736], B[736], W[735], sum[736], W[736]);
	adder a738(A[737], B[737], W[736], sum[737], W[737]);
	adder a739(A[738], B[738], W[737], sum[738], W[738]);
	adder a740(A[739], B[739], W[738], sum[739], W[739]);
	adder a741(A[740], B[740], W[739], sum[740], W[740]);
	adder a742(A[741], B[741], W[740], sum[741], W[741]);
	adder a743(A[742], B[742], W[741], sum[742], W[742]);
	adder a744(A[743], B[743], W[742], sum[743], W[743]);
	adder a745(A[744], B[744], W[743], sum[744], W[744]);
	adder a746(A[745], B[745], W[744], sum[745], W[745]);
	adder a747(A[746], B[746], W[745], sum[746], W[746]);
	adder a748(A[747], B[747], W[746], sum[747], W[747]);
	adder a749(A[748], B[748], W[747], sum[748], W[748]);
	adder a750(A[749], B[749], W[748], sum[749], W[749]);
	adder a751(A[750], B[750], W[749], sum[750], W[750]);
	adder a752(A[751], B[751], W[750], sum[751], W[751]);
	adder a753(A[752], B[752], W[751], sum[752], W[752]);
	adder a754(A[753], B[753], W[752], sum[753], W[753]);
	adder a755(A[754], B[754], W[753], sum[754], W[754]);
	adder a756(A[755], B[755], W[754], sum[755], W[755]);
	adder a757(A[756], B[756], W[755], sum[756], W[756]);
	adder a758(A[757], B[757], W[756], sum[757], W[757]);
	adder a759(A[758], B[758], W[757], sum[758], W[758]);
	adder a760(A[759], B[759], W[758], sum[759], W[759]);
	adder a761(A[760], B[760], W[759], sum[760], W[760]);
	adder a762(A[761], B[761], W[760], sum[761], W[761]);
	adder a763(A[762], B[762], W[761], sum[762], W[762]);
	adder a764(A[763], B[763], W[762], sum[763], W[763]);
	adder a765(A[764], B[764], W[763], sum[764], W[764]);
	adder a766(A[765], B[765], W[764], sum[765], W[765]);
	adder a767(A[766], B[766], W[765], sum[766], W[766]);
	adder a768(A[767], B[767], W[766], sum[767], W[767]);
	adder a769(A[768], B[768], W[767], sum[768], W[768]);
	adder a770(A[769], B[769], W[768], sum[769], W[769]);
	adder a771(A[770], B[770], W[769], sum[770], W[770]);
	adder a772(A[771], B[771], W[770], sum[771], W[771]);
	adder a773(A[772], B[772], W[771], sum[772], W[772]);
	adder a774(A[773], B[773], W[772], sum[773], W[773]);
	adder a775(A[774], B[774], W[773], sum[774], W[774]);
	adder a776(A[775], B[775], W[774], sum[775], W[775]);
	adder a777(A[776], B[776], W[775], sum[776], W[776]);
	adder a778(A[777], B[777], W[776], sum[777], W[777]);
	adder a779(A[778], B[778], W[777], sum[778], W[778]);
	adder a780(A[779], B[779], W[778], sum[779], W[779]);
	adder a781(A[780], B[780], W[779], sum[780], W[780]);
	adder a782(A[781], B[781], W[780], sum[781], W[781]);
	adder a783(A[782], B[782], W[781], sum[782], W[782]);
	adder a784(A[783], B[783], W[782], sum[783], W[783]);
	adder a785(A[784], B[784], W[783], sum[784], W[784]);
	adder a786(A[785], B[785], W[784], sum[785], W[785]);
	adder a787(A[786], B[786], W[785], sum[786], W[786]);
	adder a788(A[787], B[787], W[786], sum[787], W[787]);
	adder a789(A[788], B[788], W[787], sum[788], W[788]);
	adder a790(A[789], B[789], W[788], sum[789], W[789]);
	adder a791(A[790], B[790], W[789], sum[790], W[790]);
	adder a792(A[791], B[791], W[790], sum[791], W[791]);
	adder a793(A[792], B[792], W[791], sum[792], W[792]);
	adder a794(A[793], B[793], W[792], sum[793], W[793]);
	adder a795(A[794], B[794], W[793], sum[794], W[794]);
	adder a796(A[795], B[795], W[794], sum[795], W[795]);
	adder a797(A[796], B[796], W[795], sum[796], W[796]);
	adder a798(A[797], B[797], W[796], sum[797], W[797]);
	adder a799(A[798], B[798], W[797], sum[798], W[798]);
	adder a800(A[799], B[799], W[798], sum[799], W[799]);
	adder a801(A[800], B[800], W[799], sum[800], W[800]);
	adder a802(A[801], B[801], W[800], sum[801], W[801]);
	adder a803(A[802], B[802], W[801], sum[802], W[802]);
	adder a804(A[803], B[803], W[802], sum[803], W[803]);
	adder a805(A[804], B[804], W[803], sum[804], W[804]);
	adder a806(A[805], B[805], W[804], sum[805], W[805]);
	adder a807(A[806], B[806], W[805], sum[806], W[806]);
	adder a808(A[807], B[807], W[806], sum[807], W[807]);
	adder a809(A[808], B[808], W[807], sum[808], W[808]);
	adder a810(A[809], B[809], W[808], sum[809], W[809]);
	adder a811(A[810], B[810], W[809], sum[810], W[810]);
	adder a812(A[811], B[811], W[810], sum[811], W[811]);
	adder a813(A[812], B[812], W[811], sum[812], W[812]);
	adder a814(A[813], B[813], W[812], sum[813], W[813]);
	adder a815(A[814], B[814], W[813], sum[814], W[814]);
	adder a816(A[815], B[815], W[814], sum[815], W[815]);
	adder a817(A[816], B[816], W[815], sum[816], W[816]);
	adder a818(A[817], B[817], W[816], sum[817], W[817]);
	adder a819(A[818], B[818], W[817], sum[818], W[818]);
	adder a820(A[819], B[819], W[818], sum[819], W[819]);
	adder a821(A[820], B[820], W[819], sum[820], W[820]);
	adder a822(A[821], B[821], W[820], sum[821], W[821]);
	adder a823(A[822], B[822], W[821], sum[822], W[822]);
	adder a824(A[823], B[823], W[822], sum[823], W[823]);
	adder a825(A[824], B[824], W[823], sum[824], W[824]);
	adder a826(A[825], B[825], W[824], sum[825], W[825]);
	adder a827(A[826], B[826], W[825], sum[826], W[826]);
	adder a828(A[827], B[827], W[826], sum[827], W[827]);
	adder a829(A[828], B[828], W[827], sum[828], W[828]);
	adder a830(A[829], B[829], W[828], sum[829], W[829]);
	adder a831(A[830], B[830], W[829], sum[830], W[830]);
	adder a832(A[831], B[831], W[830], sum[831], W[831]);
	adder a833(A[832], B[832], W[831], sum[832], W[832]);
	adder a834(A[833], B[833], W[832], sum[833], W[833]);
	adder a835(A[834], B[834], W[833], sum[834], W[834]);
	adder a836(A[835], B[835], W[834], sum[835], W[835]);
	adder a837(A[836], B[836], W[835], sum[836], W[836]);
	adder a838(A[837], B[837], W[836], sum[837], W[837]);
	adder a839(A[838], B[838], W[837], sum[838], W[838]);
	adder a840(A[839], B[839], W[838], sum[839], W[839]);
	adder a841(A[840], B[840], W[839], sum[840], W[840]);
	adder a842(A[841], B[841], W[840], sum[841], W[841]);
	adder a843(A[842], B[842], W[841], sum[842], W[842]);
	adder a844(A[843], B[843], W[842], sum[843], W[843]);
	adder a845(A[844], B[844], W[843], sum[844], W[844]);
	adder a846(A[845], B[845], W[844], sum[845], W[845]);
	adder a847(A[846], B[846], W[845], sum[846], W[846]);
	adder a848(A[847], B[847], W[846], sum[847], W[847]);
	adder a849(A[848], B[848], W[847], sum[848], W[848]);
	adder a850(A[849], B[849], W[848], sum[849], W[849]);
	adder a851(A[850], B[850], W[849], sum[850], W[850]);
	adder a852(A[851], B[851], W[850], sum[851], W[851]);
	adder a853(A[852], B[852], W[851], sum[852], W[852]);
	adder a854(A[853], B[853], W[852], sum[853], W[853]);
	adder a855(A[854], B[854], W[853], sum[854], W[854]);
	adder a856(A[855], B[855], W[854], sum[855], W[855]);
	adder a857(A[856], B[856], W[855], sum[856], W[856]);
	adder a858(A[857], B[857], W[856], sum[857], W[857]);
	adder a859(A[858], B[858], W[857], sum[858], W[858]);
	adder a860(A[859], B[859], W[858], sum[859], W[859]);
	adder a861(A[860], B[860], W[859], sum[860], W[860]);
	adder a862(A[861], B[861], W[860], sum[861], W[861]);
	adder a863(A[862], B[862], W[861], sum[862], W[862]);
	adder a864(A[863], B[863], W[862], sum[863], W[863]);
	adder a865(A[864], B[864], W[863], sum[864], W[864]);
	adder a866(A[865], B[865], W[864], sum[865], W[865]);
	adder a867(A[866], B[866], W[865], sum[866], W[866]);
	adder a868(A[867], B[867], W[866], sum[867], W[867]);
	adder a869(A[868], B[868], W[867], sum[868], W[868]);
	adder a870(A[869], B[869], W[868], sum[869], W[869]);
	adder a871(A[870], B[870], W[869], sum[870], W[870]);
	adder a872(A[871], B[871], W[870], sum[871], W[871]);
	adder a873(A[872], B[872], W[871], sum[872], W[872]);
	adder a874(A[873], B[873], W[872], sum[873], W[873]);
	adder a875(A[874], B[874], W[873], sum[874], W[874]);
	adder a876(A[875], B[875], W[874], sum[875], W[875]);
	adder a877(A[876], B[876], W[875], sum[876], W[876]);
	adder a878(A[877], B[877], W[876], sum[877], W[877]);
	adder a879(A[878], B[878], W[877], sum[878], W[878]);
	adder a880(A[879], B[879], W[878], sum[879], W[879]);
	adder a881(A[880], B[880], W[879], sum[880], W[880]);
	adder a882(A[881], B[881], W[880], sum[881], W[881]);
	adder a883(A[882], B[882], W[881], sum[882], W[882]);
	adder a884(A[883], B[883], W[882], sum[883], W[883]);
	adder a885(A[884], B[884], W[883], sum[884], W[884]);
	adder a886(A[885], B[885], W[884], sum[885], W[885]);
	adder a887(A[886], B[886], W[885], sum[886], W[886]);
	adder a888(A[887], B[887], W[886], sum[887], W[887]);
	adder a889(A[888], B[888], W[887], sum[888], W[888]);
	adder a890(A[889], B[889], W[888], sum[889], W[889]);
	adder a891(A[890], B[890], W[889], sum[890], W[890]);
	adder a892(A[891], B[891], W[890], sum[891], W[891]);
	adder a893(A[892], B[892], W[891], sum[892], W[892]);
	adder a894(A[893], B[893], W[892], sum[893], W[893]);
	adder a895(A[894], B[894], W[893], sum[894], W[894]);
	adder a896(A[895], B[895], W[894], sum[895], W[895]);
	adder a897(A[896], B[896], W[895], sum[896], W[896]);
	adder a898(A[897], B[897], W[896], sum[897], W[897]);
	adder a899(A[898], B[898], W[897], sum[898], W[898]);
	adder a900(A[899], B[899], W[898], sum[899], W[899]);
	adder a901(A[900], B[900], W[899], sum[900], W[900]);
	adder a902(A[901], B[901], W[900], sum[901], W[901]);
	adder a903(A[902], B[902], W[901], sum[902], W[902]);
	adder a904(A[903], B[903], W[902], sum[903], W[903]);
	adder a905(A[904], B[904], W[903], sum[904], W[904]);
	adder a906(A[905], B[905], W[904], sum[905], W[905]);
	adder a907(A[906], B[906], W[905], sum[906], W[906]);
	adder a908(A[907], B[907], W[906], sum[907], W[907]);
	adder a909(A[908], B[908], W[907], sum[908], W[908]);
	adder a910(A[909], B[909], W[908], sum[909], W[909]);
	adder a911(A[910], B[910], W[909], sum[910], W[910]);
	adder a912(A[911], B[911], W[910], sum[911], W[911]);
	adder a913(A[912], B[912], W[911], sum[912], W[912]);
	adder a914(A[913], B[913], W[912], sum[913], W[913]);
	adder a915(A[914], B[914], W[913], sum[914], W[914]);
	adder a916(A[915], B[915], W[914], sum[915], W[915]);
	adder a917(A[916], B[916], W[915], sum[916], W[916]);
	adder a918(A[917], B[917], W[916], sum[917], W[917]);
	adder a919(A[918], B[918], W[917], sum[918], W[918]);
	adder a920(A[919], B[919], W[918], sum[919], W[919]);
	adder a921(A[920], B[920], W[919], sum[920], W[920]);
	adder a922(A[921], B[921], W[920], sum[921], W[921]);
	adder a923(A[922], B[922], W[921], sum[922], W[922]);
	adder a924(A[923], B[923], W[922], sum[923], W[923]);
	adder a925(A[924], B[924], W[923], sum[924], W[924]);
	adder a926(A[925], B[925], W[924], sum[925], W[925]);
	adder a927(A[926], B[926], W[925], sum[926], W[926]);
	adder a928(A[927], B[927], W[926], sum[927], W[927]);
	adder a929(A[928], B[928], W[927], sum[928], W[928]);
	adder a930(A[929], B[929], W[928], sum[929], W[929]);
	adder a931(A[930], B[930], W[929], sum[930], W[930]);
	adder a932(A[931], B[931], W[930], sum[931], W[931]);
	adder a933(A[932], B[932], W[931], sum[932], W[932]);
	adder a934(A[933], B[933], W[932], sum[933], W[933]);
	adder a935(A[934], B[934], W[933], sum[934], W[934]);
	adder a936(A[935], B[935], W[934], sum[935], W[935]);
	adder a937(A[936], B[936], W[935], sum[936], W[936]);
	adder a938(A[937], B[937], W[936], sum[937], W[937]);
	adder a939(A[938], B[938], W[937], sum[938], W[938]);
	adder a940(A[939], B[939], W[938], sum[939], W[939]);
	adder a941(A[940], B[940], W[939], sum[940], W[940]);
	adder a942(A[941], B[941], W[940], sum[941], W[941]);
	adder a943(A[942], B[942], W[941], sum[942], W[942]);
	adder a944(A[943], B[943], W[942], sum[943], W[943]);
	adder a945(A[944], B[944], W[943], sum[944], W[944]);
	adder a946(A[945], B[945], W[944], sum[945], W[945]);
	adder a947(A[946], B[946], W[945], sum[946], W[946]);
	adder a948(A[947], B[947], W[946], sum[947], W[947]);
	adder a949(A[948], B[948], W[947], sum[948], W[948]);
	adder a950(A[949], B[949], W[948], sum[949], W[949]);
	adder a951(A[950], B[950], W[949], sum[950], W[950]);
	adder a952(A[951], B[951], W[950], sum[951], W[951]);
	adder a953(A[952], B[952], W[951], sum[952], W[952]);
	adder a954(A[953], B[953], W[952], sum[953], W[953]);
	adder a955(A[954], B[954], W[953], sum[954], W[954]);
	adder a956(A[955], B[955], W[954], sum[955], W[955]);
	adder a957(A[956], B[956], W[955], sum[956], W[956]);
	adder a958(A[957], B[957], W[956], sum[957], W[957]);
	adder a959(A[958], B[958], W[957], sum[958], W[958]);
	adder a960(A[959], B[959], W[958], sum[959], W[959]);
	adder a961(A[960], B[960], W[959], sum[960], W[960]);
	adder a962(A[961], B[961], W[960], sum[961], W[961]);
	adder a963(A[962], B[962], W[961], sum[962], W[962]);
	adder a964(A[963], B[963], W[962], sum[963], W[963]);
	adder a965(A[964], B[964], W[963], sum[964], W[964]);
	adder a966(A[965], B[965], W[964], sum[965], W[965]);
	adder a967(A[966], B[966], W[965], sum[966], W[966]);
	adder a968(A[967], B[967], W[966], sum[967], W[967]);
	adder a969(A[968], B[968], W[967], sum[968], W[968]);
	adder a970(A[969], B[969], W[968], sum[969], W[969]);
	adder a971(A[970], B[970], W[969], sum[970], W[970]);
	adder a972(A[971], B[971], W[970], sum[971], W[971]);
	adder a973(A[972], B[972], W[971], sum[972], W[972]);
	adder a974(A[973], B[973], W[972], sum[973], W[973]);
	adder a975(A[974], B[974], W[973], sum[974], W[974]);
	adder a976(A[975], B[975], W[974], sum[975], W[975]);
	adder a977(A[976], B[976], W[975], sum[976], W[976]);
	adder a978(A[977], B[977], W[976], sum[977], W[977]);
	adder a979(A[978], B[978], W[977], sum[978], W[978]);
	adder a980(A[979], B[979], W[978], sum[979], W[979]);
	adder a981(A[980], B[980], W[979], sum[980], W[980]);
	adder a982(A[981], B[981], W[980], sum[981], W[981]);
	adder a983(A[982], B[982], W[981], sum[982], W[982]);
	adder a984(A[983], B[983], W[982], sum[983], W[983]);
	adder a985(A[984], B[984], W[983], sum[984], W[984]);
	adder a986(A[985], B[985], W[984], sum[985], W[985]);
	adder a987(A[986], B[986], W[985], sum[986], W[986]);
	adder a988(A[987], B[987], W[986], sum[987], W[987]);
	adder a989(A[988], B[988], W[987], sum[988], W[988]);
	adder a990(A[989], B[989], W[988], sum[989], W[989]);
	adder a991(A[990], B[990], W[989], sum[990], W[990]);
	adder a992(A[991], B[991], W[990], sum[991], W[991]);
	adder a993(A[992], B[992], W[991], sum[992], W[992]);
	adder a994(A[993], B[993], W[992], sum[993], W[993]);
	adder a995(A[994], B[994], W[993], sum[994], W[994]);
	adder a996(A[995], B[995], W[994], sum[995], W[995]);
	adder a997(A[996], B[996], W[995], sum[996], W[996]);
	adder a998(A[997], B[997], W[996], sum[997], W[997]);
	adder a999(A[998], B[998], W[997], sum[998], W[998]);
	adder a1000(A[999], B[999], W[998], sum[999], W[999]);
	adder a1001(A[1000], B[1000], W[999], sum[1000], W[1000]);
	adder a1002(A[1001], B[1001], W[1000], sum[1001], W[1001]);
	adder a1003(A[1002], B[1002], W[1001], sum[1002], W[1002]);
	adder a1004(A[1003], B[1003], W[1002], sum[1003], W[1003]);
	adder a1005(A[1004], B[1004], W[1003], sum[1004], W[1004]);
	adder a1006(A[1005], B[1005], W[1004], sum[1005], W[1005]);
	adder a1007(A[1006], B[1006], W[1005], sum[1006], W[1006]);
	adder a1008(A[1007], B[1007], W[1006], sum[1007], W[1007]);
	adder a1009(A[1008], B[1008], W[1007], sum[1008], W[1008]);
	adder a1010(A[1009], B[1009], W[1008], sum[1009], W[1009]);
	adder a1011(A[1010], B[1010], W[1009], sum[1010], W[1010]);
	adder a1012(A[1011], B[1011], W[1010], sum[1011], W[1011]);
	adder a1013(A[1012], B[1012], W[1011], sum[1012], W[1012]);
	adder a1014(A[1013], B[1013], W[1012], sum[1013], W[1013]);
	adder a1015(A[1014], B[1014], W[1013], sum[1014], W[1014]);
	adder a1016(A[1015], B[1015], W[1014], sum[1015], W[1015]);
	adder a1017(A[1016], B[1016], W[1015], sum[1016], W[1016]);
	adder a1018(A[1017], B[1017], W[1016], sum[1017], W[1017]);
	adder a1019(A[1018], B[1018], W[1017], sum[1018], W[1018]);
	adder a1020(A[1019], B[1019], W[1018], sum[1019], W[1019]);
	adder a1021(A[1020], B[1020], W[1019], sum[1020], W[1020]);
	adder a1022(A[1021], B[1021], W[1020], sum[1021], W[1021]);
	adder a1023(A[1022], B[1022], W[1021], sum[1022], W[1022]);
	adder a1024(A[1023], B[1023], W[1022], sum[1023], W[1023]);

	assign Cout = W[1023];

endmodule