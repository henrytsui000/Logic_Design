module check_zero(A, Q);
	input [1023:0] A;
	output Q;
	wire ret;

	or ans(ret, A[1023], A[1022], A[1021], A[1020], A[1019], A[1018], A[1017], A[1016], A[1015], A[1014], A[1013], A[1012], A[1011], A[1010], A[1009], A[1008], A[1007], A[1006], A[1005], A[1004], A[1003], A[1002], A[1001], A[1000], A[999], A[998], A[997], A[996], A[995], A[994], A[993], A[992], A[991], A[990], A[989], A[988], A[987], A[986], A[985], A[984], A[983], A[982], A[981], A[980], A[979], A[978], A[977], A[976], A[975], A[974], A[973], A[972], A[971], A[970], A[969], A[968], A[967], A[966], A[965], A[964], A[963], A[962], A[961], A[960], A[959], A[958], A[957], A[956], A[955], A[954], A[953], A[952], A[951], A[950], A[949], A[948], A[947], A[946], A[945], A[944], A[943], A[942], A[941], A[940], A[939], A[938], A[937], A[936], A[935], A[934], A[933], A[932], A[931], A[930], A[929], A[928], A[927], A[926], A[925], A[924], A[923], A[922], A[921], A[920], A[919], A[918], A[917], A[916], A[915], A[914], A[913], A[912], A[911], A[910], A[909], A[908], A[907], A[906], A[905], A[904], A[903], A[902], A[901], A[900], A[899], A[898], A[897], A[896], A[895], A[894], A[893], A[892], A[891], A[890], A[889], A[888], A[887], A[886], A[885], A[884], A[883], A[882], A[881], A[880], A[879], A[878], A[877], A[876], A[875], A[874], A[873], A[872], A[871], A[870], A[869], A[868], A[867], A[866], A[865], A[864], A[863], A[862], A[861], A[860], A[859], A[858], A[857], A[856], A[855], A[854], A[853], A[852], A[851], A[850], A[849], A[848], A[847], A[846], A[845], A[844], A[843], A[842], A[841], A[840], A[839], A[838], A[837], A[836], A[835], A[834], A[833], A[832], A[831], A[830], A[829], A[828], A[827], A[826], A[825], A[824], A[823], A[822], A[821], A[820], A[819], A[818], A[817], A[816], A[815], A[814], A[813], A[812], A[811], A[810], A[809], A[808], A[807], A[806], A[805], A[804], A[803], A[802], A[801], A[800], A[799], A[798], A[797], A[796], A[795], A[794], A[793], A[792], A[791], A[790], A[789], A[788], A[787], A[786], A[785], A[784], A[783], A[782], A[781], A[780], A[779], A[778], A[777], A[776], A[775], A[774], A[773], A[772], A[771], A[770], A[769], A[768], A[767], A[766], A[765], A[764], A[763], A[762], A[761], A[760], A[759], A[758], A[757], A[756], A[755], A[754], A[753], A[752], A[751], A[750], A[749], A[748], A[747], A[746], A[745], A[744], A[743], A[742], A[741], A[740], A[739], A[738], A[737], A[736], A[735], A[734], A[733], A[732], A[731], A[730], A[729], A[728], A[727], A[726], A[725], A[724], A[723], A[722], A[721], A[720], A[719], A[718], A[717], A[716], A[715], A[714], A[713], A[712], A[711], A[710], A[709], A[708], A[707], A[706], A[705], A[704], A[703], A[702], A[701], A[700], A[699], A[698], A[697], A[696], A[695], A[694], A[693], A[692], A[691], A[690], A[689], A[688], A[687], A[686], A[685], A[684], A[683], A[682], A[681], A[680], A[679], A[678], A[677], A[676], A[675], A[674], A[673], A[672], A[671], A[670], A[669], A[668], A[667], A[666], A[665], A[664], A[663], A[662], A[661], A[660], A[659], A[658], A[657], A[656], A[655], A[654], A[653], A[652], A[651], A[650], A[649], A[648], A[647], A[646], A[645], A[644], A[643], A[642], A[641], A[640], A[639], A[638], A[637], A[636], A[635], A[634], A[633], A[632], A[631], A[630], A[629], A[628], A[627], A[626], A[625], A[624], A[623], A[622], A[621], A[620], A[619], A[618], A[617], A[616], A[615], A[614], A[613], A[612], A[611], A[610], A[609], A[608], A[607], A[606], A[605], A[604], A[603], A[602], A[601], A[600], A[599], A[598], A[597], A[596], A[595], A[594], A[593], A[592], A[591], A[590], A[589], A[588], A[587], A[586], A[585], A[584], A[583], A[582], A[581], A[580], A[579], A[578], A[577], A[576], A[575], A[574], A[573], A[572], A[571], A[570], A[569], A[568], A[567], A[566], A[565], A[564], A[563], A[562], A[561], A[560], A[559], A[558], A[557], A[556], A[555], A[554], A[553], A[552], A[551], A[550], A[549], A[548], A[547], A[546], A[545], A[544], A[543], A[542], A[541], A[540], A[539], A[538], A[537], A[536], A[535], A[534], A[533], A[532], A[531], A[530], A[529], A[528], A[527], A[526], A[525], A[524], A[523], A[522], A[521], A[520], A[519], A[518], A[517], A[516], A[515], A[514], A[513], A[512], A[511], A[510], A[509], A[508], A[507], A[506], A[505], A[504], A[503], A[502], A[501], A[500], A[499], A[498], A[497], A[496], A[495], A[494], A[493], A[492], A[491], A[490], A[489], A[488], A[487], A[486], A[485], A[484], A[483], A[482], A[481], A[480], A[479], A[478], A[477], A[476], A[475], A[474], A[473], A[472], A[471], A[470], A[469], A[468], A[467], A[466], A[465], A[464], A[463], A[462], A[461], A[460], A[459], A[458], A[457], A[456], A[455], A[454], A[453], A[452], A[451], A[450], A[449], A[448], A[447], A[446], A[445], A[444], A[443], A[442], A[441], A[440], A[439], A[438], A[437], A[436], A[435], A[434], A[433], A[432], A[431], A[430], A[429], A[428], A[427], A[426], A[425], A[424], A[423], A[422], A[421], A[420], A[419], A[418], A[417], A[416], A[415], A[414], A[413], A[412], A[411], A[410], A[409], A[408], A[407], A[406], A[405], A[404], A[403], A[402], A[401], A[400], A[399], A[398], A[397], A[396], A[395], A[394], A[393], A[392], A[391], A[390], A[389], A[388], A[387], A[386], A[385], A[384], A[383], A[382], A[381], A[380], A[379], A[378], A[377], A[376], A[375], A[374], A[373], A[372], A[371], A[370], A[369], A[368], A[367], A[366], A[365], A[364], A[363], A[362], A[361], A[360], A[359], A[358], A[357], A[356], A[355], A[354], A[353], A[352], A[351], A[350], A[349], A[348], A[347], A[346], A[345], A[344], A[343], A[342], A[341], A[340], A[339], A[338], A[337], A[336], A[335], A[334], A[333], A[332], A[331], A[330], A[329], A[328], A[327], A[326], A[325], A[324], A[323], A[322], A[321], A[320], A[319], A[318], A[317], A[316], A[315], A[314], A[313], A[312], A[311], A[310], A[309], A[308], A[307], A[306], A[305], A[304], A[303], A[302], A[301], A[300], A[299], A[298], A[297], A[296], A[295], A[294], A[293], A[292], A[291], A[290], A[289], A[288], A[287], A[286], A[285], A[284], A[283], A[282], A[281], A[280], A[279], A[278], A[277], A[276], A[275], A[274], A[273], A[272], A[271], A[270], A[269], A[268], A[267], A[266], A[265], A[264], A[263], A[262], A[261], A[260], A[259], A[258], A[257], A[256], A[255], A[254], A[253], A[252], A[251], A[250], A[249], A[248], A[247], A[246], A[245], A[244], A[243], A[242], A[241], A[240], A[239], A[238], A[237], A[236], A[235], A[234], A[233], A[232], A[231], A[230], A[229], A[228], A[227], A[226], A[225], A[224], A[223], A[222], A[221], A[220], A[219], A[218], A[217], A[216], A[215], A[214], A[213], A[212], A[211], A[210], A[209], A[208], A[207], A[206], A[205], A[204], A[203], A[202], A[201], A[200], A[199], A[198], A[197], A[196], A[195], A[194], A[193], A[192], A[191], A[190], A[189], A[188], A[187], A[186], A[185], A[184], A[183], A[182], A[181], A[180], A[179], A[178], A[177], A[176], A[175], A[174], A[173], A[172], A[171], A[170], A[169], A[168], A[167], A[166], A[165], A[164], A[163], A[162], A[161], A[160], A[159], A[158], A[157], A[156], A[155], A[154], A[153], A[152], A[151], A[150], A[149], A[148], A[147], A[146], A[145], A[144], A[143], A[142], A[141], A[140], A[139], A[138], A[137], A[136], A[135], A[134], A[133], A[132], A[131], A[130], A[129], A[128], A[127], A[126], A[125], A[124], A[123], A[122], A[121], A[120], A[119], A[118], A[117], A[116], A[115], A[114], A[113], A[112], A[111], A[110], A[109], A[108], A[107], A[106], A[105], A[104], A[103], A[102], A[101], A[100], A[99], A[98], A[97], A[96], A[95], A[94], A[93], A[92], A[91], A[90], A[89], A[88], A[87], A[86], A[85], A[84], A[83], A[82], A[81], A[80], A[79], A[78], A[77], A[76], A[75], A[74], A[73], A[72], A[71], A[70], A[69], A[68], A[67], A[66], A[65], A[64], A[63], A[62], A[61], A[60], A[59], A[58], A[57], A[56], A[55], A[54], A[53], A[52], A[51], A[50], A[49], A[48], A[47], A[46], A[45], A[44], A[43], A[42], A[41], A[40], A[39], A[38], A[37], A[36], A[35], A[34], A[33], A[32], A[31], A[30], A[29], A[28], A[27], A[26], A[25], A[24], A[23], A[22], A[21], A[20], A[19], A[18], A[17], A[16], A[15], A[14], A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], A[5], A[4], A[3], A[2], A[1], A[0]);
	not not1(Q, ret);
endmodule